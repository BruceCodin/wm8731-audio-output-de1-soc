// pll.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module pll (
		input  wire        clk_clk,                           //                     clk.clk
		output wire        clock_12_clk,                      //                clock_12.clk
		input  wire        onchip_memory2_0_reset1_reset,     // onchip_memory2_0_reset1.reset
		input  wire        onchip_memory2_0_reset1_reset_req, //                        .reset_req
		input  wire [17:0] onchip_memory2_0_s1_address,       //     onchip_memory2_0_s1.address
		input  wire        onchip_memory2_0_s1_debugaccess,   //                        .debugaccess
		input  wire        onchip_memory2_0_s1_clken,         //                        .clken
		input  wire        onchip_memory2_0_s1_chipselect,    //                        .chipselect
		input  wire        onchip_memory2_0_s1_write,         //                        .write
		output wire [15:0] onchip_memory2_0_s1_readdata,      //                        .readdata
		input  wire [15:0] onchip_memory2_0_s1_writedata,     //                        .writedata
		input  wire [1:0]  onchip_memory2_0_s1_byteenable,    //                        .byteenable
		input  wire        reset_reset_n                      //                   reset.reset_n
	);

	wire    pll_0_outclk1_clk; // pll_0:outclk_1 -> onchip_memory2_0:clk

	pll_onchip_memory2_0 onchip_memory2_0 (
		.clk         (pll_0_outclk1_clk),                 //   clk1.clk
		.address     (onchip_memory2_0_s1_address),       //     s1.address
		.debugaccess (onchip_memory2_0_s1_debugaccess),   //       .debugaccess
		.clken       (onchip_memory2_0_s1_clken),         //       .clken
		.chipselect  (onchip_memory2_0_s1_chipselect),    //       .chipselect
		.write       (onchip_memory2_0_s1_write),         //       .write
		.readdata    (onchip_memory2_0_s1_readdata),      //       .readdata
		.writedata   (onchip_memory2_0_s1_writedata),     //       .writedata
		.byteenable  (onchip_memory2_0_s1_byteenable),    //       .byteenable
		.reset       (onchip_memory2_0_reset1_reset),     // reset1.reset
		.reset_req   (onchip_memory2_0_reset1_reset_req), //       .reset_req
		.freeze      (1'b0)                               // (terminated)
	);

	pll_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (clock_12_clk),      // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   // (terminated)
	);

endmodule
